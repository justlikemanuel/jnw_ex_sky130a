magic
tech sky130A
magscale 1 2
timestamp 1736461524
<< locali >>
rect -106 -368 86 168
rect 1046 -368 1238 170
rect -106 -372 1370 -368
rect -106 -552 284 -372
rect 464 -552 1370 -372
rect -106 -560 1370 -552
<< viali >>
rect 284 -552 464 -372
<< metal1 >>
rect 986 3946 1036 4231
rect 146 2293 210 3868
rect 658 3754 1036 3946
rect 140 2227 146 2293
rect 212 2227 218 2293
rect 146 104 210 2227
rect 275 443 465 3589
rect 986 3137 1036 3754
rect 763 3087 1036 3137
rect 717 2293 783 2299
rect 717 2221 783 2227
rect 986 1479 1036 3087
rect 771 1429 1036 1479
rect 986 653 1036 1429
rect 773 603 1036 653
rect 278 -372 470 320
rect 986 42 1036 603
rect 278 -552 284 -372
rect 464 -552 470 -372
rect 278 -564 470 -552
<< via1 >>
rect 146 2227 212 2293
rect 717 2227 783 2293
<< metal2 >>
rect 146 2293 212 2299
rect 212 2227 717 2293
rect 783 2227 789 2293
rect 146 2221 212 2227
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1736460924
transform 1 0 -14 0 1 3214
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1736460924
transform 1 0 -10 0 1 16
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1736460924
transform 1 0 -12 0 1 814
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1736460924
transform 1 0 -12 0 1 1614
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1736460924
transform 1 0 -12 0 1 2414
box -184 -128 1336 928
<< labels >>
flabel metal2 212 2227 717 2293 0 FreeSans 1600 0 0 0 IBPS_5U
port 1 nsew
flabel locali 464 -560 1370 -368 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel metal1 658 3754 1036 3946 0 FreeSans 1600 0 0 0 IBNS_20U
port 3 nsew
<< end >>
